-------------------------------------------------------------------------------
-- Projeto: Projeto Genius
-- Curso: Engenharia de Sistemas Turma PN5
--
-- Integrantes:
--   Guilherme Fachinelli
--   Rafael Campello Soares
--   Gustavo Silvestre Barroso
--
-- Descrição:
--   Arquivo pertencente ao projeto digital baseado no jogo Genius.
--   Desenvolvido para fins acadêmicos na disciplina de Sistemas Digitais.
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.all;

entity tb_Sequence_design is
end tb_Sequence_design;

architecture sim of tb_Sequence_design is

    function slv_to_string(slv: std_logic_vector) return string is
        variable result : string(1 to slv'length);
    begin
        for i in slv'range loop
            case slv(i) is
                when '0' => result(i - slv'low + 1) := '0';
                when '1' => result(i - slv'low + 1) := '1';
                when 'U' => result(i - slv'low + 1) := 'U';
                when 'X' => result(i - slv'low + 1) := 'X';
                when 'Z' => result(i - slv'low + 1) := 'Z';
                when others => result(i - slv'low + 1) := '?';
            end case;
        end loop;
        return result;
    end function;

    constant CLK_PERIOD : time := 10 ns;

    signal clk      : std_logic := '0';
    signal rst      : std_logic := '0';
    signal start    : std_logic := '0';
    signal base_out : array_3X7bits;
    signal done     : std_logic;

begin

    -- UUT ----------------------------------------------------
    uut: entity work.Sequence_design
        port map (
            clk       => clk,
            rst       => rst,
            start     => start,
            base_out  => base_out,
            ready_out => done
        );

    -- Clock ---------------------------------------------------
    clk_process : process
    begin
        report "[CLK] Clock process iniciado" severity note;
        while true loop
            clk <= '0'; wait for CLK_PERIOD/2;
            clk <= '1'; wait for CLK_PERIOD/2;
        end loop;
    end process;

    -- Estímulos 
    stim_proc : process
    begin
        report "[TB] Testbench iniciado" severity note;

        -- Reset
        rst <= '1';
        report "[TB] Reset = 1" severity note;
        wait for 30 ns;

        rst <= '0';
        report "[TB] Reset = 0" severity note;

        wait for 721 ns;

        -- Start
        start <= '1';
        report "[TB] Start = 1" severity note;
        wait for CLK_PERIOD;
        start <= '0';
        report "[TB] Start = 0" severity note;

        wait for 100 ns;

        report "[TB] Esperando done..." severity note;

        wait until done = '1' for 100000 ns;

        if done = '1' then
            report "[TB] DONE = 1 RECEBIDO" severity note;

            report "=== Resultado base_out ===";
            for i in base_out'range loop
                report "base_out(" & integer'image(i) & ") = " &
                       slv_to_string(base_out(i)) & " (" &
                       integer'image(to_integer(unsigned(base_out(i)))) & ")";
            end loop;

        else
            report "ERRO: Módulo não completou dentro do tempo esperado!" severity error;
        end if;

        report "=== Simulação encerrada ===";
        assert false report "STOP" severity failure;
        wait;

    end process;

end sim;
